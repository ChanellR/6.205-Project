  module particle_buffer(
    input wire clk_in, 
    input wire rst_in, 
    input wire busy, 
    output logic [47:0] p_out, 
    output logic p_valid_out
  );

  logic [$clog2(200)-1:0] addr;

  logic [200:0][47:0] buffer = {48'h4411c5484444,
48'h43773c1fc33b,
48'hc0394374c294,
48'h2f85be19c5cd,
48'h408dc29c4222,
48'h339c45843b5d,
48'hbcc6457fc52e,
48'hc4b441434495,
48'hc05ec0b0443a,
48'hc572b9d5c572,
48'hc4153eccc181,
48'h44b63e8fbd2a,
48'hc0693a62bba6,
48'h3c973961c175,
48'hbef53cae44b2,
48'h4496bfb243ef,
48'hc43bc21fbc2c,
48'h44a8c58cc58d,
48'h4164402ec1c5,
48'h45bf4551c39c,
48'hc47bc460c484,
48'hc17cbc454128,
48'hbba440b83fc3,
48'hbc424421c5cf,
48'h450d3a2ec1d4,
48'hc4753f534098,
48'h44bf4015c2ed,
48'h4248c4e6c457,
48'h4029c38243ca,
48'hb58d37ba3d06,
48'h401bc5ccc2b5,
48'hc457451cc459,
48'hb971c1b0be86,
48'h4415bf964490,
48'hc5c94565c471,
48'hc1ed43834437,
48'hc56dc44f3e38,
48'h45754517c54d,
48'h440d4440442f,
48'hc547b91bc111,
48'hc22745823784,
48'h423a3d074592,
48'hc448c08abaac,
48'h44bf43fec537,
48'hc2c43af7c1d7,
48'h3bd4bd15b682,
48'h3fe4c3fc42d3,
48'h410a45bb440c,
48'h40e1bdf3c280,
48'hc5c540fcb95a,
48'hc301c2c7b7ca,
48'hbec14534411b,
48'h446ac1be440d,
48'h4481c4d7bcc5,
48'h3f66453940d2,
48'hb840bf634286,
48'hb2c5c4994497,
48'h4407c43dc155,
48'h44784457c52b,
48'hb683c15c44b5,
48'hc2633db74147,
48'h3b5fbd4bc527,
48'h3c3e3208c06b,
48'hb11bc4cd4045,
48'h3782c4e7c4c1,
48'h4020c330c2f9,
48'h42dfb7e3b41f,
48'hc189bf634367,
48'hc5fa441e41cc,
48'h417c4190c5a4,
48'hc25dc222c54b,
48'hc5f9c1edbd54,
48'hc2c13556c46f,
48'hc36a406bc58a,
48'hc36f3f94c4c1,
48'hc0e3c4c4c4eb,
48'hc5f5bc01c04a,
48'h41dbc2623d2e,
48'h44aa3f07b5c0,
48'h41eec255c529,
48'hb57243c1bd39,
48'h40703e38c326,
48'h30f73f44431e,
48'h3ea52c43c5b1,
48'hc5f7c2403342,
48'h2dcfc31f444d,
48'h3843c501c40c,
48'hb846c446ba33,
48'hc48443d942f9,
48'h32724551c4a1,
48'h45393f00c372,
48'hbbe043584172,
48'hbeb7b8183fdb,
48'haec5369e3f7c,
48'h3e21c5e03d18,
48'hc36cbc94bccf,
48'hc1cec1ccc52f,
48'h43dd45c5bcda,
48'h43d8458f4330,
48'hc4cebfe6c2e2,
48'hbbb7c57543a6,
48'h3ccc258cbf0a,
48'hc4ef414cc387,
48'hb9b4432ec4ab,
48'hb989c3e439fc,
48'hbfd23d844168,
48'h432ec44a3d8b,
48'h420242a244a1,
48'hc509412944ab,
48'hbc6d44404207,
48'hc26842a843f7,
48'h3e4340ccc506,
48'h3ebdc1aa33b1,
48'hbc7d3976c513,
48'h44abb7f1c4e2,
48'h43ec40e84421,
48'hc1453d29c4e5,
48'h3ece3d37c07e,
48'hbcb5c36ebc51,
48'h45fe3e4f3f2a,
48'h41d7c394c35a,
48'hc1d437d945ca,
48'h3947c05d437b,
48'hc53642473e00,
48'hc1ba430345e9,
48'hc5df4083c090,
48'hb65141e1c0ba,
48'h4391bc314403,
48'h45944434c4b7,
48'h457744764083,
48'h45e6458cb62e,
48'hc35145584310,
48'h3d1ac2ed45ec,
48'h456ebf9a3a6b,
48'h43f4b98a4156,
48'hc4cf455a43b9,
48'h3c213f734342,
48'h3fbd41f8c238,
48'hc5a1c025422d,
48'hc325c4f9456e,
48'h3b363d15c562,
48'h44f4c075b97c,
48'hc23eba7d45c7,
48'h442f40f745f8,
48'h40f83eb0bc09,
48'h36b8c1c03046,
48'hc22eb6fe3f17,
48'hc53041b6c4c4,
48'hb73fc0d94485,
48'h3d5ec5fbb540,
48'h369d3ed043fd,
48'hc20fc4f2b6d2,
48'hc5b2c2e3c34d,
48'ha8e440a040f6,
48'hc4b8bedc40fe,
48'hbe04c463c52c,
48'h45c04525c004,
48'h445444f1bc86,
48'h3f0b37e13f09,
48'h449ec4953c6b,
48'hc0724475c2bf,
48'h3d9cb5c63cf7,
48'hb9ee3a48b452,
48'h3773b8f844c8,
48'hc4bd417c4253,
48'hc440c275c53a,
48'hc5e3441fc433,
48'hb097c015c433,
48'hc59b38b64009,
48'h4420c5ad4595,
48'h38e3c4eac47e,
48'h3ed8b06d420a,
48'hc022bcbab032,
48'hc36840b7c056,
48'h3e6c40eebf8d,
48'hc1e044d24588,
48'hbed23d323c3f,
48'h445ec0f9b92f,
48'h2f8ec1073295,
48'h44a340e1be51,
48'h3e034131b5ba,
48'h443742034513,
48'h4400c25a4266,
48'hc347c58140b4,
48'h42b4442445ad,
48'h446fc4ec3834,
48'h3e46c30ac27e,
48'hc042c557b00b,
48'hc4ffb4583a04,
48'h4508c4bb3f76,
48'h403d437a4599,
48'h3c0442efc529,
48'h4455c38ac355,
48'hc22fc5a4b8ac,
48'hc4df427e43d9,
48'h4000be93406a,
48'hc5a3c4574429,
48'hc587c0ef45e6,
48'h3a44c328bf37,
48'h40e3bba74599}; 

  // xilinx_true_dual_port_read_first_2_clock_ram #(
  //   .RAM_WIDTH(48),                       // Specify RAM data width
  //   .RAM_DEPTH(200),                     // Specify RAM depth (number of entries)
  //   .RAM_PERFORMANCE("HIGH_PERFORMANCE"), // Select "HIGH_PERFORMANCE" or "LOW_LATENCY"
  //   .INIT_FILE("../../data/pb.mem")                        // Specify name/location of RAM initialization file if using one (leave blank if not)
  // ) your_instance_name (
  //   .addra(addr),   // Port A address bus, width determined from RAM_DEPTH
  //   .addrb(),   // Port B address bus, width determined from RAM_DEPTH
  //   .dina(),     // Port A RAM input data, width determined from RAM_WIDTH
  //   .dinb(),     // Port B RAM input data, width determined from RAM_WIDTH
  //   .clka(clk_in),     // Port A clock
  //   .clkb(clk_in),     // Port B clock
  //   .wea(1'b0),       // Port A write enable
  //   .web(1'b0),       // Port B write enable
  //   .ena(1'b1),       // Port A RAM Enable, for additional power savings, disable port when not in use
  //   .enb(1'b1),       // Port B RAM Enable, for additional power savings, disable port when not in use
  //   .rsta(rst_in),     // Port A output reset (does not affect memory contents)
  //   .rstb(rst_in),     // Port B output reset (does not affect memory contents)
  //   .regcea(1'b1), // Port A output register enable
  //   .regceb(1'b1), // Port B output register enable
  //   .douta(),   // Port A RAM output data, width determined from RAM_WIDTH
  //   .doutb(p_out)    // Port B RAM output data, width determined from RAM_WIDTH
  // );

  always_ff @(posedge clk_in) begin
    if(rst_in) begin 
      addr <=0; 
    end else begin 
      if(~busy) begin 
        addr <= addr + 1;
        p_valid_out <= 1;  
        p_out <= buffer[addr]; 
      end else begin 
        p_valid_out <= 0; 
      end
    end
  end 

endmodule 
