//    tmds_encoder tmds_red(
//        .clk_in(clk_pixel),
//        .rst_in(sys_rst_pixel),
//        .data_in(red),
//        .control_in(2'b0),
//        .ve_in(ad_pipe),
//        .tmds_out(tmds_10b[2]));

//    tmds_encoder tmds_green(
//          .clk_in(clk_pixel),
//          .rst_in(sys_rst_pixel),
//          .data_in(green),
//          .control_in(2'b0),
//          .ve_in(ad_pipe),
//          .tmds_out(tmds_10b[1]));

//    tmds_encoder tmds_blue(
//         .clk_in(clk_pixel),
//         .rst_in(sys_rst_pixel),
//         .data_in(blue),
//         .control_in({vsync_pipe,hsync_pipe}),
//         .ve_in(ad_pipe),
//         .tmds_out(tmds_10b[0]));

  
//    //three tmds_serializers (blue, green, red):
//    //MISSING: two more serializers for the green and blue tmds signals.
//    tmds_serializer red_ser(
//          .clk_pixel_in(clk_pixel),
//          .clk_5x_in(clk_5x),
//          .rst_in(sys_rst_pixel),
//          .tmds_in(tmds_10b[2]),
//          .tmds_out(tmds_signal[2]));
//    tmds_serializer green_ser(
//          .clk_pixel_in(clk_pixel),
//          .clk_5x_in(clk_5x),
//          .rst_in(sys_rst_pixel),
//          .tmds_in(tmds_10b[1]),
//          .tmds_out(tmds_signal[1]));
//    tmds_serializer blue_ser(
//          .clk_pixel_in(clk_pixel),
//          .clk_5x_in(clk_5x),
//          .rst_in(sys_rst_pixel),
//          .tmds_in(tmds_10b[0]),
//          .tmds_out(tmds_signal[0]));

//    //output buffers generating differential signals:
//    //three for the r,g,b signals and one that is at the pixel clock rate
//    //the HDMI receivers use recover logic coupled with the control signals asserted
//    //during blanking and sync periods to synchronize their faster bit clocks off
//    //of the slower pixel clock (so they can recover a clock of about 742.5 MHz from
//    //the slower 74.25 MHz clock)
//    OBUFDS OBUFDS_blue (.I(tmds_signal[0]), .O(hdmi_tx_p[0]), .OB(hdmi_tx_n[0]));
//    OBUFDS OBUFDS_green(.I(tmds_signal[1]), .O(hdmi_tx_p[1]), .OB(hdmi_tx_n[1]));
//    OBUFDS OBUFDS_red  (.I(tmds_signal[2]), .O(hdmi_tx_p[2]), .OB(hdmi_tx_n[2]));
//    OBUFDS OBUFDS_clock(.I(clk_pixel), .O(hdmi_clk_p), .OB(hdmi_clk_n));